// qsys_fpga_emif.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module qsys_fpga_emif (
		input  wire         clk_clk,                                       //                          clk.clk
		input  wire         emif_fm_0_local_reset_req_local_reset_req,     //    emif_fm_0_local_reset_req.local_reset_req
		output wire         emif_fm_0_local_reset_status_local_reset_done, // emif_fm_0_local_reset_status.local_reset_done
		input  wire         emif_fm_0_oct_oct_rzqin,                       //                emif_fm_0_oct.oct_rzqin
		output wire [0:0]   emif_fm_0_mem_mem_ck,                          //                emif_fm_0_mem.mem_ck
		output wire [0:0]   emif_fm_0_mem_mem_ck_n,                        //                             .mem_ck_n
		output wire [16:0]  emif_fm_0_mem_mem_a,                           //                             .mem_a
		output wire [0:0]   emif_fm_0_mem_mem_act_n,                       //                             .mem_act_n
		output wire [1:0]   emif_fm_0_mem_mem_ba,                          //                             .mem_ba
		output wire [0:0]   emif_fm_0_mem_mem_bg,                          //                             .mem_bg
		output wire [0:0]   emif_fm_0_mem_mem_cke,                         //                             .mem_cke
		output wire [0:0]   emif_fm_0_mem_mem_cs_n,                        //                             .mem_cs_n
		output wire [0:0]   emif_fm_0_mem_mem_odt,                         //                             .mem_odt
		output wire [0:0]   emif_fm_0_mem_mem_reset_n,                     //                             .mem_reset_n
		output wire [0:0]   emif_fm_0_mem_mem_par,                         //                             .mem_par
		input  wire [0:0]   emif_fm_0_mem_mem_alert_n,                     //                             .mem_alert_n
		inout  wire [1:0]   emif_fm_0_mem_mem_dqs,                         //                             .mem_dqs
		inout  wire [1:0]   emif_fm_0_mem_mem_dqs_n,                       //                             .mem_dqs_n
		inout  wire [15:0]  emif_fm_0_mem_mem_dq,                          //                             .mem_dq
		inout  wire [1:0]   emif_fm_0_mem_mem_dbi_n,                       //                             .mem_dbi_n
		output wire         emif_fm_0_status_local_cal_success,            //             emif_fm_0_status.local_cal_success
		output wire         emif_fm_0_status_local_cal_fail,               //                             .local_cal_fail
		output wire         emif_fm_0_emif_usr_reset_n_reset_n,            //   emif_fm_0_emif_usr_reset_n.reset_n
		output wire         emif_fm_0_emif_usr_clk_clk,                    //       emif_fm_0_emif_usr_clk.clk
		output wire         emif_fm_0_ctrl_amm_0_waitrequest_n,            //         emif_fm_0_ctrl_amm_0.waitrequest_n
		input  wire         emif_fm_0_ctrl_amm_0_read,                     //                             .read
		input  wire         emif_fm_0_ctrl_amm_0_write,                    //                             .write
		input  wire [26:0]  emif_fm_0_ctrl_amm_0_address,                  //                             .address
		output wire [127:0] emif_fm_0_ctrl_amm_0_readdata,                 //                             .readdata
		input  wire [127:0] emif_fm_0_ctrl_amm_0_writedata,                //                             .writedata
		input  wire [6:0]   emif_fm_0_ctrl_amm_0_burstcount,               //                             .burstcount
		input  wire [15:0]  emif_fm_0_ctrl_amm_0_byteenable,               //                             .byteenable
		output wire         emif_fm_0_ctrl_amm_0_readdatavalid,            //                             .readdatavalid
		input  wire         reset_reset_n                                  //                        reset.reset_n
	);

	wire           emif_cal_0_emif_calbus_clk_clk;             // emif_cal_0:calbus_clk -> emif_fm_0:calbus_clk
	wire           clock_in_out_clk_clk;                       // clock_in:out_clk -> [emif_cal_0:cal_debug_clk_clk, emif_fm_0:pll_ref_clk, reset_in:clk]
	wire    [31:0] emif_cal_0_emif_calbus_0_calbus_wdata;      // emif_cal_0:calbus_wdata_0 -> emif_fm_0:calbus_wdata
	wire    [19:0] emif_cal_0_emif_calbus_0_calbus_address;    // emif_cal_0:calbus_address_0 -> emif_fm_0:calbus_address
	wire  [4095:0] emif_fm_0_emif_calbus_calbus_seq_param_tbl; // emif_fm_0:calbus_seq_param_tbl -> emif_cal_0:calbus_seq_param_tbl_0
	wire           emif_cal_0_emif_calbus_0_calbus_read;       // emif_cal_0:calbus_read_0 -> emif_fm_0:calbus_read
	wire           emif_cal_0_emif_calbus_0_calbus_write;      // emif_cal_0:calbus_write_0 -> emif_fm_0:calbus_write
	wire    [31:0] emif_fm_0_emif_calbus_calbus_rdata;         // emif_fm_0:calbus_rdata -> emif_cal_0:calbus_rdata_0
	wire           reset_in_out_reset_reset;                   // reset_in:out_reset_n -> emif_cal_0:cal_debug_reset_n_reset

	qsys_fpga_emif_clock_in clock_in (
		.in_clk  (clk_clk),              //   input,  width = 1,  in_clk.clk
		.out_clk (clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	qsys_fpga_emif_emif_cal_0 emif_cal_0 (
		.calbus_read_0           (emif_cal_0_emif_calbus_0_calbus_read),       //  output,     width = 1,     emif_calbus_0.calbus_read
		.calbus_write_0          (emif_cal_0_emif_calbus_0_calbus_write),      //  output,     width = 1,                  .calbus_write
		.calbus_address_0        (emif_cal_0_emif_calbus_0_calbus_address),    //  output,    width = 20,                  .calbus_address
		.calbus_wdata_0          (emif_cal_0_emif_calbus_0_calbus_wdata),      //  output,    width = 32,                  .calbus_wdata
		.calbus_rdata_0          (emif_fm_0_emif_calbus_calbus_rdata),         //   input,    width = 32,                  .calbus_rdata
		.calbus_seq_param_tbl_0  (emif_fm_0_emif_calbus_calbus_seq_param_tbl), //   input,  width = 4096,                  .calbus_seq_param_tbl
		.calbus_clk              (emif_cal_0_emif_calbus_clk_clk),             //  output,     width = 1,   emif_calbus_clk.clk
		.cal_debug_clk_clk       (clock_in_out_clk_clk),                       //   input,     width = 1,     cal_debug_clk.clk
		.cal_debug_reset_n_reset (~reset_in_out_reset_reset)                   //   input,     width = 1, cal_debug_reset_n.reset
	);

	qsys_fpga_emif_emif_fm_0 emif_fm_0 (
		.local_reset_req      (emif_fm_0_local_reset_req_local_reset_req),     //   input,     width = 1,    local_reset_req.local_reset_req
		.local_reset_done     (emif_fm_0_local_reset_status_local_reset_done), //  output,     width = 1, local_reset_status.local_reset_done
		.pll_ref_clk          (clock_in_out_clk_clk),                          //   input,     width = 1,        pll_ref_clk.clk
		.oct_rzqin            (emif_fm_0_oct_oct_rzqin),                       //   input,     width = 1,                oct.oct_rzqin
		.mem_ck               (emif_fm_0_mem_mem_ck),                          //  output,     width = 1,                mem.mem_ck
		.mem_ck_n             (emif_fm_0_mem_mem_ck_n),                        //  output,     width = 1,                   .mem_ck_n
		.mem_a                (emif_fm_0_mem_mem_a),                           //  output,    width = 17,                   .mem_a
		.mem_act_n            (emif_fm_0_mem_mem_act_n),                       //  output,     width = 1,                   .mem_act_n
		.mem_ba               (emif_fm_0_mem_mem_ba),                          //  output,     width = 2,                   .mem_ba
		.mem_bg               (emif_fm_0_mem_mem_bg),                          //  output,     width = 1,                   .mem_bg
		.mem_cke              (emif_fm_0_mem_mem_cke),                         //  output,     width = 1,                   .mem_cke
		.mem_cs_n             (emif_fm_0_mem_mem_cs_n),                        //  output,     width = 1,                   .mem_cs_n
		.mem_odt              (emif_fm_0_mem_mem_odt),                         //  output,     width = 1,                   .mem_odt
		.mem_reset_n          (emif_fm_0_mem_mem_reset_n),                     //  output,     width = 1,                   .mem_reset_n
		.mem_par              (emif_fm_0_mem_mem_par),                         //  output,     width = 1,                   .mem_par
		.mem_alert_n          (emif_fm_0_mem_mem_alert_n),                     //   input,     width = 1,                   .mem_alert_n
		.mem_dqs              (emif_fm_0_mem_mem_dqs),                         //   inout,     width = 2,                   .mem_dqs
		.mem_dqs_n            (emif_fm_0_mem_mem_dqs_n),                       //   inout,     width = 2,                   .mem_dqs_n
		.mem_dq               (emif_fm_0_mem_mem_dq),                          //   inout,    width = 16,                   .mem_dq
		.mem_dbi_n            (emif_fm_0_mem_mem_dbi_n),                       //   inout,     width = 2,                   .mem_dbi_n
		.local_cal_success    (emif_fm_0_status_local_cal_success),            //  output,     width = 1,             status.local_cal_success
		.local_cal_fail       (emif_fm_0_status_local_cal_fail),               //  output,     width = 1,                   .local_cal_fail
		.emif_usr_reset_n     (emif_fm_0_emif_usr_reset_n_reset_n),            //  output,     width = 1,   emif_usr_reset_n.reset_n
		.emif_usr_clk         (emif_fm_0_emif_usr_clk_clk),                    //  output,     width = 1,       emif_usr_clk.clk
		.amm_ready_0          (emif_fm_0_ctrl_amm_0_waitrequest_n),            //  output,     width = 1,         ctrl_amm_0.waitrequest_n
		.amm_read_0           (emif_fm_0_ctrl_amm_0_read),                     //   input,     width = 1,                   .read
		.amm_write_0          (emif_fm_0_ctrl_amm_0_write),                    //   input,     width = 1,                   .write
		.amm_address_0        (emif_fm_0_ctrl_amm_0_address),                  //   input,    width = 27,                   .address
		.amm_readdata_0       (emif_fm_0_ctrl_amm_0_readdata),                 //  output,   width = 128,                   .readdata
		.amm_writedata_0      (emif_fm_0_ctrl_amm_0_writedata),                //   input,   width = 128,                   .writedata
		.amm_burstcount_0     (emif_fm_0_ctrl_amm_0_burstcount),               //   input,     width = 7,                   .burstcount
		.amm_byteenable_0     (emif_fm_0_ctrl_amm_0_byteenable),               //   input,    width = 16,                   .byteenable
		.amm_readdatavalid_0  (emif_fm_0_ctrl_amm_0_readdatavalid),            //  output,     width = 1,                   .readdatavalid
		.calbus_read          (emif_cal_0_emif_calbus_0_calbus_read),          //   input,     width = 1,        emif_calbus.calbus_read
		.calbus_write         (emif_cal_0_emif_calbus_0_calbus_write),         //   input,     width = 1,                   .calbus_write
		.calbus_address       (emif_cal_0_emif_calbus_0_calbus_address),       //   input,    width = 20,                   .calbus_address
		.calbus_wdata         (emif_cal_0_emif_calbus_0_calbus_wdata),         //   input,    width = 32,                   .calbus_wdata
		.calbus_rdata         (emif_fm_0_emif_calbus_calbus_rdata),            //  output,    width = 32,                   .calbus_rdata
		.calbus_seq_param_tbl (emif_fm_0_emif_calbus_calbus_seq_param_tbl),    //  output,  width = 4096,                   .calbus_seq_param_tbl
		.calbus_clk           (emif_cal_0_emif_calbus_clk_clk)                 //   input,     width = 1,    emif_calbus_clk.clk
	);

	qsys_fpga_emif_reset_in reset_in (
		.clk         (clock_in_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_reset_n),            //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_in_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

endmodule
